module XOR(
    input a,b,
    output c
);
  
  assign c = a ^ b ;

endmodule